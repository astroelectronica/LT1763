.title KiCad schematic
.include "C:/AE/LT1763/_models/C3216X5R2A105K160AA_s.mod"
.include "C:/AE/LT1763/_models/CEU4J2X7R2A103K125AE_s.mod"
.include "C:/AE/LT1763/_models/CGA5L3X5R1H106K160AB_s.mod"
.include "C:/AE/LT1763/_models/LT1763.lib"
R2 /VOUT /ADJ {RADJU}
XU3 /BYP /VOUT CEU4J2X7R2A103K125AE_s
R3 /ADJ 0 {RADJB}
I1 /VOUT 0 {ILOAD}
XU4 /VOUT 0 CGA5L3X5R1H106K160AB_s
V1 /VIN 0 {VSOURCE}
XU1 /VIN 0 C3216X5R2A105K160AA_s
XU2 /VOUT /ADJ 0 /BYP /VIN /VIN LT1763
.end
